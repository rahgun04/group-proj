// unsaved.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module unsaved (
		output wire [31:0] atan2_a_external_connection_export,      //      atan2_a_external_connection.export
		output wire [31:0] atan2_b_external_connection_export,      //      atan2_b_external_connection.export
		input  wire [31:0] atan2_q_external_connection_export,      //      atan2_q_external_connection.export
		input  wire        clk_clk,                                 //                              clk.clk
		input  wire        i2c_busy_external_connection_export,     //     i2c_busy_external_connection.export
		output wire [7:0]  i2c_dev_addr_external_connection_export, // i2c_dev_addr_external_connection.export
		output wire        i2c_en_external_connection_export,       //       i2c_en_external_connection.export
		input  wire [7:0]  i2c_miso_external_connection_export,     //     i2c_miso_external_connection.export
		output wire [7:0]  i2c_mosi_external_connection_export,     //     i2c_mosi_external_connection.export
		output wire [7:0]  i2c_reg_addr_external_connection_export, // i2c_reg_addr_external_connection.export
		output wire        i2c_rst_external_connection_export,      //      i2c_rst_external_connection.export
		output wire        i2c_rw_external_connection_export,       //       i2c_rw_external_connection.export
		input  wire [31:0] in_l_external_connection_export,         //         in_l_external_connection.export
		output wire [9:0]  led_external_connection_export,          //          led_external_connection.export
		output wire [31:0] out0_external_connection_export,         //         out0_external_connection.export
		output wire [31:0] out1_external_connection_export,         //         out1_external_connection.export
		input  wire        reset_reset_n,                           //                            reset.reset_n
		output wire        sample_clk_external_connection_export    //   sample_clk_external_connection.export
	);

	wire  [31:0] cpu_data_master_readdata;                                  // mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	wire         cpu_data_master_waitrequest;                               // mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	wire         cpu_data_master_debugaccess;                               // cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	wire  [17:0] cpu_data_master_address;                                   // cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	wire   [3:0] cpu_data_master_byteenable;                                // cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	wire         cpu_data_master_read;                                      // cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	wire         cpu_data_master_write;                                     // cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	wire  [31:0] cpu_data_master_writedata;                                 // cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	wire  [31:0] cpu_instruction_master_readdata;                           // mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	wire         cpu_instruction_master_waitrequest;                        // mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	wire  [17:0] cpu_instruction_master_address;                            // cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	wire         cpu_instruction_master_read;                               // cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;    // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest; // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_readdata;            // cpu:debug_mem_slave_readdata -> mm_interconnect_0:cpu_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu_debug_mem_slave_waitrequest;         // cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu_debug_mem_slave_debugaccess;         // mm_interconnect_0:cpu_debug_mem_slave_debugaccess -> cpu:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_debug_mem_slave_address;             // mm_interconnect_0:cpu_debug_mem_slave_address -> cpu:debug_mem_slave_address
	wire         mm_interconnect_0_cpu_debug_mem_slave_read;                // mm_interconnect_0:cpu_debug_mem_slave_read -> cpu:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu_debug_mem_slave_byteenable;          // mm_interconnect_0:cpu_debug_mem_slave_byteenable -> cpu:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu_debug_mem_slave_write;               // mm_interconnect_0:cpu_debug_mem_slave_write -> cpu:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_writedata;           // mm_interconnect_0:cpu_debug_mem_slave_writedata -> cpu:debug_mem_slave_writedata
	wire         mm_interconnect_0_led_s1_chipselect;                       // mm_interconnect_0:led_s1_chipselect -> led:chipselect
	wire  [31:0] mm_interconnect_0_led_s1_readdata;                         // led:readdata -> mm_interconnect_0:led_s1_readdata
	wire   [1:0] mm_interconnect_0_led_s1_address;                          // mm_interconnect_0:led_s1_address -> led:address
	wire         mm_interconnect_0_led_s1_write;                            // mm_interconnect_0:led_s1_write -> led:write_n
	wire  [31:0] mm_interconnect_0_led_s1_writedata;                        // mm_interconnect_0:led_s1_writedata -> led:writedata
	wire         mm_interconnect_0_onchip_memory_s1_chipselect;             // mm_interconnect_0:onchip_memory_s1_chipselect -> onchip_memory:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory_s1_readdata;               // onchip_memory:readdata -> mm_interconnect_0:onchip_memory_s1_readdata
	wire  [13:0] mm_interconnect_0_onchip_memory_s1_address;                // mm_interconnect_0:onchip_memory_s1_address -> onchip_memory:address
	wire   [3:0] mm_interconnect_0_onchip_memory_s1_byteenable;             // mm_interconnect_0:onchip_memory_s1_byteenable -> onchip_memory:byteenable
	wire         mm_interconnect_0_onchip_memory_s1_write;                  // mm_interconnect_0:onchip_memory_s1_write -> onchip_memory:write
	wire  [31:0] mm_interconnect_0_onchip_memory_s1_writedata;              // mm_interconnect_0:onchip_memory_s1_writedata -> onchip_memory:writedata
	wire         mm_interconnect_0_onchip_memory_s1_clken;                  // mm_interconnect_0:onchip_memory_s1_clken -> onchip_memory:clken
	wire         mm_interconnect_0_out0_s1_chipselect;                      // mm_interconnect_0:out0_s1_chipselect -> out0:chipselect
	wire  [31:0] mm_interconnect_0_out0_s1_readdata;                        // out0:readdata -> mm_interconnect_0:out0_s1_readdata
	wire   [1:0] mm_interconnect_0_out0_s1_address;                         // mm_interconnect_0:out0_s1_address -> out0:address
	wire         mm_interconnect_0_out0_s1_write;                           // mm_interconnect_0:out0_s1_write -> out0:write_n
	wire  [31:0] mm_interconnect_0_out0_s1_writedata;                       // mm_interconnect_0:out0_s1_writedata -> out0:writedata
	wire         mm_interconnect_0_out1_s1_chipselect;                      // mm_interconnect_0:out1_s1_chipselect -> out1:chipselect
	wire  [31:0] mm_interconnect_0_out1_s1_readdata;                        // out1:readdata -> mm_interconnect_0:out1_s1_readdata
	wire   [1:0] mm_interconnect_0_out1_s1_address;                         // mm_interconnect_0:out1_s1_address -> out1:address
	wire         mm_interconnect_0_out1_s1_write;                           // mm_interconnect_0:out1_s1_write -> out1:write_n
	wire  [31:0] mm_interconnect_0_out1_s1_writedata;                       // mm_interconnect_0:out1_s1_writedata -> out1:writedata
	wire  [31:0] mm_interconnect_0_in_h_s1_readdata;                        // in_H:readdata -> mm_interconnect_0:in_H_s1_readdata
	wire   [1:0] mm_interconnect_0_in_h_s1_address;                         // mm_interconnect_0:in_H_s1_address -> in_H:address
	wire  [31:0] mm_interconnect_0_in_l_s1_readdata;                        // in_L:readdata -> mm_interconnect_0:in_L_s1_readdata
	wire   [1:0] mm_interconnect_0_in_l_s1_address;                         // mm_interconnect_0:in_L_s1_address -> in_L:address
	wire         mm_interconnect_0_sample_clk_s1_chipselect;                // mm_interconnect_0:sample_clk_s1_chipselect -> sample_clk:chipselect
	wire  [31:0] mm_interconnect_0_sample_clk_s1_readdata;                  // sample_clk:readdata -> mm_interconnect_0:sample_clk_s1_readdata
	wire   [1:0] mm_interconnect_0_sample_clk_s1_address;                   // mm_interconnect_0:sample_clk_s1_address -> sample_clk:address
	wire         mm_interconnect_0_sample_clk_s1_write;                     // mm_interconnect_0:sample_clk_s1_write -> sample_clk:write_n
	wire  [31:0] mm_interconnect_0_sample_clk_s1_writedata;                 // mm_interconnect_0:sample_clk_s1_writedata -> sample_clk:writedata
	wire         mm_interconnect_0_i2c_rst_s1_chipselect;                   // mm_interconnect_0:i2c_rst_s1_chipselect -> i2c_rst:chipselect
	wire  [31:0] mm_interconnect_0_i2c_rst_s1_readdata;                     // i2c_rst:readdata -> mm_interconnect_0:i2c_rst_s1_readdata
	wire   [1:0] mm_interconnect_0_i2c_rst_s1_address;                      // mm_interconnect_0:i2c_rst_s1_address -> i2c_rst:address
	wire         mm_interconnect_0_i2c_rst_s1_write;                        // mm_interconnect_0:i2c_rst_s1_write -> i2c_rst:write_n
	wire  [31:0] mm_interconnect_0_i2c_rst_s1_writedata;                    // mm_interconnect_0:i2c_rst_s1_writedata -> i2c_rst:writedata
	wire         mm_interconnect_0_i2c_en_s1_chipselect;                    // mm_interconnect_0:i2c_en_s1_chipselect -> i2c_en:chipselect
	wire  [31:0] mm_interconnect_0_i2c_en_s1_readdata;                      // i2c_en:readdata -> mm_interconnect_0:i2c_en_s1_readdata
	wire   [1:0] mm_interconnect_0_i2c_en_s1_address;                       // mm_interconnect_0:i2c_en_s1_address -> i2c_en:address
	wire         mm_interconnect_0_i2c_en_s1_write;                         // mm_interconnect_0:i2c_en_s1_write -> i2c_en:write_n
	wire  [31:0] mm_interconnect_0_i2c_en_s1_writedata;                     // mm_interconnect_0:i2c_en_s1_writedata -> i2c_en:writedata
	wire         mm_interconnect_0_i2c_rw_s1_chipselect;                    // mm_interconnect_0:i2c_rw_s1_chipselect -> i2c_rw:chipselect
	wire  [31:0] mm_interconnect_0_i2c_rw_s1_readdata;                      // i2c_rw:readdata -> mm_interconnect_0:i2c_rw_s1_readdata
	wire   [1:0] mm_interconnect_0_i2c_rw_s1_address;                       // mm_interconnect_0:i2c_rw_s1_address -> i2c_rw:address
	wire         mm_interconnect_0_i2c_rw_s1_write;                         // mm_interconnect_0:i2c_rw_s1_write -> i2c_rw:write_n
	wire  [31:0] mm_interconnect_0_i2c_rw_s1_writedata;                     // mm_interconnect_0:i2c_rw_s1_writedata -> i2c_rw:writedata
	wire         mm_interconnect_0_i2c_mosi_s1_chipselect;                  // mm_interconnect_0:i2c_mosi_s1_chipselect -> i2c_mosi:chipselect
	wire  [31:0] mm_interconnect_0_i2c_mosi_s1_readdata;                    // i2c_mosi:readdata -> mm_interconnect_0:i2c_mosi_s1_readdata
	wire   [1:0] mm_interconnect_0_i2c_mosi_s1_address;                     // mm_interconnect_0:i2c_mosi_s1_address -> i2c_mosi:address
	wire         mm_interconnect_0_i2c_mosi_s1_write;                       // mm_interconnect_0:i2c_mosi_s1_write -> i2c_mosi:write_n
	wire  [31:0] mm_interconnect_0_i2c_mosi_s1_writedata;                   // mm_interconnect_0:i2c_mosi_s1_writedata -> i2c_mosi:writedata
	wire         mm_interconnect_0_i2c_reg_addr_s1_chipselect;              // mm_interconnect_0:i2c_reg_addr_s1_chipselect -> i2c_reg_addr:chipselect
	wire  [31:0] mm_interconnect_0_i2c_reg_addr_s1_readdata;                // i2c_reg_addr:readdata -> mm_interconnect_0:i2c_reg_addr_s1_readdata
	wire   [1:0] mm_interconnect_0_i2c_reg_addr_s1_address;                 // mm_interconnect_0:i2c_reg_addr_s1_address -> i2c_reg_addr:address
	wire         mm_interconnect_0_i2c_reg_addr_s1_write;                   // mm_interconnect_0:i2c_reg_addr_s1_write -> i2c_reg_addr:write_n
	wire  [31:0] mm_interconnect_0_i2c_reg_addr_s1_writedata;               // mm_interconnect_0:i2c_reg_addr_s1_writedata -> i2c_reg_addr:writedata
	wire         mm_interconnect_0_i2c_dev_addr_s1_chipselect;              // mm_interconnect_0:i2c_dev_addr_s1_chipselect -> i2c_dev_addr:chipselect
	wire  [31:0] mm_interconnect_0_i2c_dev_addr_s1_readdata;                // i2c_dev_addr:readdata -> mm_interconnect_0:i2c_dev_addr_s1_readdata
	wire   [1:0] mm_interconnect_0_i2c_dev_addr_s1_address;                 // mm_interconnect_0:i2c_dev_addr_s1_address -> i2c_dev_addr:address
	wire         mm_interconnect_0_i2c_dev_addr_s1_write;                   // mm_interconnect_0:i2c_dev_addr_s1_write -> i2c_dev_addr:write_n
	wire  [31:0] mm_interconnect_0_i2c_dev_addr_s1_writedata;               // mm_interconnect_0:i2c_dev_addr_s1_writedata -> i2c_dev_addr:writedata
	wire  [31:0] mm_interconnect_0_i2c_miso_s1_readdata;                    // i2c_miso:readdata -> mm_interconnect_0:i2c_miso_s1_readdata
	wire   [1:0] mm_interconnect_0_i2c_miso_s1_address;                     // mm_interconnect_0:i2c_miso_s1_address -> i2c_miso:address
	wire  [31:0] mm_interconnect_0_i2c_busy_s1_readdata;                    // i2c_busy:readdata -> mm_interconnect_0:i2c_busy_s1_readdata
	wire   [1:0] mm_interconnect_0_i2c_busy_s1_address;                     // mm_interconnect_0:i2c_busy_s1_address -> i2c_busy:address
	wire         mm_interconnect_0_atan2_a_s1_chipselect;                   // mm_interconnect_0:atan2_a_s1_chipselect -> atan2_a:chipselect
	wire  [31:0] mm_interconnect_0_atan2_a_s1_readdata;                     // atan2_a:readdata -> mm_interconnect_0:atan2_a_s1_readdata
	wire   [1:0] mm_interconnect_0_atan2_a_s1_address;                      // mm_interconnect_0:atan2_a_s1_address -> atan2_a:address
	wire         mm_interconnect_0_atan2_a_s1_write;                        // mm_interconnect_0:atan2_a_s1_write -> atan2_a:write_n
	wire  [31:0] mm_interconnect_0_atan2_a_s1_writedata;                    // mm_interconnect_0:atan2_a_s1_writedata -> atan2_a:writedata
	wire         mm_interconnect_0_atan2_b_s1_chipselect;                   // mm_interconnect_0:atan2_b_s1_chipselect -> atan2_b:chipselect
	wire  [31:0] mm_interconnect_0_atan2_b_s1_readdata;                     // atan2_b:readdata -> mm_interconnect_0:atan2_b_s1_readdata
	wire   [1:0] mm_interconnect_0_atan2_b_s1_address;                      // mm_interconnect_0:atan2_b_s1_address -> atan2_b:address
	wire         mm_interconnect_0_atan2_b_s1_write;                        // mm_interconnect_0:atan2_b_s1_write -> atan2_b:write_n
	wire  [31:0] mm_interconnect_0_atan2_b_s1_writedata;                    // mm_interconnect_0:atan2_b_s1_writedata -> atan2_b:writedata
	wire  [31:0] mm_interconnect_0_atan2_q_s1_readdata;                     // atan2_q:readdata -> mm_interconnect_0:atan2_q_s1_readdata
	wire   [1:0] mm_interconnect_0_atan2_q_s1_address;                      // mm_interconnect_0:atan2_q_s1_address -> atan2_q:address
	wire         irq_mapper_receiver0_irq;                                  // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] cpu_irq_irq;                                               // irq_mapper:sender_irq -> cpu:irq
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [atan2_a:reset_n, atan2_b:reset_n, atan2_q:reset_n, cpu:reset_n, i2c_busy:reset_n, i2c_dev_addr:reset_n, i2c_en:reset_n, i2c_miso:reset_n, i2c_mosi:reset_n, i2c_reg_addr:reset_n, i2c_rst:reset_n, i2c_rw:reset_n, in_H:reset_n, in_L:reset_n, irq_mapper:reset, jtag_uart:rst_n, led:reset_n, mm_interconnect_0:cpu_reset_reset_bridge_in_reset_reset, onchip_memory:reset, out0:reset_n, out1:reset_n, rst_translator:in_reset, sample_clk:reset_n]
	wire         rst_controller_reset_out_reset_req;                        // rst_controller:reset_req -> [cpu:reset_req, onchip_memory:reset_req, rst_translator:reset_req_in]

	unsaved_atan2_a atan2_a (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_atan2_a_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_atan2_a_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_atan2_a_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_atan2_a_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_atan2_a_s1_readdata),   //                    .readdata
		.out_port   (atan2_a_external_connection_export)       // external_connection.export
	);

	unsaved_atan2_a atan2_b (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_atan2_b_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_atan2_b_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_atan2_b_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_atan2_b_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_atan2_b_s1_readdata),   //                    .readdata
		.out_port   (atan2_b_external_connection_export)       // external_connection.export
	);

	unsaved_atan2_q atan2_q (
		.clk      (clk_clk),                               //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address  (mm_interconnect_0_atan2_q_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_atan2_q_s1_readdata), //                    .readdata
		.in_port  (atan2_q_external_connection_export)     // external_connection.export
	);

	unsaved_cpu cpu (
		.clk                                 (clk_clk),                                           //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                   //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                //                          .reset_req
		.d_address                           (cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_data_master_read),                              //                          .read
		.d_readdata                          (cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_data_master_write),                             //                          .write
		.d_writedata                         (cpu_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                  //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                   // custom_instruction_master.readra
	);

	unsaved_i2c_busy i2c_busy (
		.clk      (clk_clk),                                //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address  (mm_interconnect_0_i2c_busy_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_i2c_busy_s1_readdata), //                    .readdata
		.in_port  (i2c_busy_external_connection_export)     // external_connection.export
	);

	unsaved_i2c_dev_addr i2c_dev_addr (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_i2c_dev_addr_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_i2c_dev_addr_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_i2c_dev_addr_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_i2c_dev_addr_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_i2c_dev_addr_s1_readdata),   //                    .readdata
		.out_port   (i2c_dev_addr_external_connection_export)       // external_connection.export
	);

	unsaved_i2c_en i2c_en (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_i2c_en_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_i2c_en_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_i2c_en_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_i2c_en_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_i2c_en_s1_readdata),   //                    .readdata
		.out_port   (i2c_en_external_connection_export)       // external_connection.export
	);

	unsaved_i2c_miso i2c_miso (
		.clk      (clk_clk),                                //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address  (mm_interconnect_0_i2c_miso_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_i2c_miso_s1_readdata), //                    .readdata
		.in_port  (i2c_miso_external_connection_export)     // external_connection.export
	);

	unsaved_i2c_dev_addr i2c_mosi (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_i2c_mosi_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_i2c_mosi_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_i2c_mosi_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_i2c_mosi_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_i2c_mosi_s1_readdata),   //                    .readdata
		.out_port   (i2c_mosi_external_connection_export)       // external_connection.export
	);

	unsaved_i2c_dev_addr i2c_reg_addr (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_i2c_reg_addr_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_i2c_reg_addr_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_i2c_reg_addr_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_i2c_reg_addr_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_i2c_reg_addr_s1_readdata),   //                    .readdata
		.out_port   (i2c_reg_addr_external_connection_export)       // external_connection.export
	);

	unsaved_i2c_en i2c_rst (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_i2c_rst_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_i2c_rst_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_i2c_rst_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_i2c_rst_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_i2c_rst_s1_readdata),   //                    .readdata
		.out_port   (i2c_rst_external_connection_export)       // external_connection.export
	);

	unsaved_i2c_en i2c_rw (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_i2c_rw_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_i2c_rw_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_i2c_rw_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_i2c_rw_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_i2c_rw_s1_readdata),   //                    .readdata
		.out_port   (i2c_rw_external_connection_export)       // external_connection.export
	);

	unsaved_atan2_q in_h (
		.clk      (clk_clk),                            //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),    //               reset.reset_n
		.address  (mm_interconnect_0_in_h_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_in_h_s1_readdata), //                    .readdata
		.in_port  ()                                    // external_connection.export
	);

	unsaved_atan2_q in_l (
		.clk      (clk_clk),                            //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),    //               reset.reset_n
		.address  (mm_interconnect_0_in_l_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_in_l_s1_readdata), //                    .readdata
		.in_port  (in_l_external_connection_export)     // external_connection.export
	);

	unsaved_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	unsaved_led led (
		.clk        (clk_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led_s1_readdata),   //                    .readdata
		.out_port   (led_external_connection_export)       // external_connection.export
	);

	unsaved_onchip_memory onchip_memory (
		.clk        (clk_clk),                                       //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),            //       .reset_req
		.freeze     (1'b0)                                           // (terminated)
	);

	unsaved_atan2_a out0 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_out0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_out0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_out0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_out0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_out0_s1_readdata),   //                    .readdata
		.out_port   (out0_external_connection_export)       // external_connection.export
	);

	unsaved_atan2_a out1 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_out1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_out1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_out1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_out1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_out1_s1_readdata),   //                    .readdata
		.out_port   (out1_external_connection_export)       // external_connection.export
	);

	unsaved_i2c_en sample_clk (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_sample_clk_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sample_clk_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sample_clk_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sample_clk_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sample_clk_s1_readdata),   //                    .readdata
		.out_port   (sample_clk_external_connection_export)       // external_connection.export
	);

	unsaved_mm_interconnect_0 mm_interconnect_0 (
		.clk_clk_clk                             (clk_clk),                                                   //                         clk_clk.clk
		.cpu_reset_reset_bridge_in_reset_reset   (rst_controller_reset_out_reset),                            // cpu_reset_reset_bridge_in_reset.reset
		.cpu_data_master_address                 (cpu_data_master_address),                                   //                 cpu_data_master.address
		.cpu_data_master_waitrequest             (cpu_data_master_waitrequest),                               //                                .waitrequest
		.cpu_data_master_byteenable              (cpu_data_master_byteenable),                                //                                .byteenable
		.cpu_data_master_read                    (cpu_data_master_read),                                      //                                .read
		.cpu_data_master_readdata                (cpu_data_master_readdata),                                  //                                .readdata
		.cpu_data_master_write                   (cpu_data_master_write),                                     //                                .write
		.cpu_data_master_writedata               (cpu_data_master_writedata),                                 //                                .writedata
		.cpu_data_master_debugaccess             (cpu_data_master_debugaccess),                               //                                .debugaccess
		.cpu_instruction_master_address          (cpu_instruction_master_address),                            //          cpu_instruction_master.address
		.cpu_instruction_master_waitrequest      (cpu_instruction_master_waitrequest),                        //                                .waitrequest
		.cpu_instruction_master_read             (cpu_instruction_master_read),                               //                                .read
		.cpu_instruction_master_readdata         (cpu_instruction_master_readdata),                           //                                .readdata
		.atan2_a_s1_address                      (mm_interconnect_0_atan2_a_s1_address),                      //                      atan2_a_s1.address
		.atan2_a_s1_write                        (mm_interconnect_0_atan2_a_s1_write),                        //                                .write
		.atan2_a_s1_readdata                     (mm_interconnect_0_atan2_a_s1_readdata),                     //                                .readdata
		.atan2_a_s1_writedata                    (mm_interconnect_0_atan2_a_s1_writedata),                    //                                .writedata
		.atan2_a_s1_chipselect                   (mm_interconnect_0_atan2_a_s1_chipselect),                   //                                .chipselect
		.atan2_b_s1_address                      (mm_interconnect_0_atan2_b_s1_address),                      //                      atan2_b_s1.address
		.atan2_b_s1_write                        (mm_interconnect_0_atan2_b_s1_write),                        //                                .write
		.atan2_b_s1_readdata                     (mm_interconnect_0_atan2_b_s1_readdata),                     //                                .readdata
		.atan2_b_s1_writedata                    (mm_interconnect_0_atan2_b_s1_writedata),                    //                                .writedata
		.atan2_b_s1_chipselect                   (mm_interconnect_0_atan2_b_s1_chipselect),                   //                                .chipselect
		.atan2_q_s1_address                      (mm_interconnect_0_atan2_q_s1_address),                      //                      atan2_q_s1.address
		.atan2_q_s1_readdata                     (mm_interconnect_0_atan2_q_s1_readdata),                     //                                .readdata
		.cpu_debug_mem_slave_address             (mm_interconnect_0_cpu_debug_mem_slave_address),             //             cpu_debug_mem_slave.address
		.cpu_debug_mem_slave_write               (mm_interconnect_0_cpu_debug_mem_slave_write),               //                                .write
		.cpu_debug_mem_slave_read                (mm_interconnect_0_cpu_debug_mem_slave_read),                //                                .read
		.cpu_debug_mem_slave_readdata            (mm_interconnect_0_cpu_debug_mem_slave_readdata),            //                                .readdata
		.cpu_debug_mem_slave_writedata           (mm_interconnect_0_cpu_debug_mem_slave_writedata),           //                                .writedata
		.cpu_debug_mem_slave_byteenable          (mm_interconnect_0_cpu_debug_mem_slave_byteenable),          //                                .byteenable
		.cpu_debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_debug_mem_slave_waitrequest),         //                                .waitrequest
		.cpu_debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_debug_mem_slave_debugaccess),         //                                .debugaccess
		.i2c_busy_s1_address                     (mm_interconnect_0_i2c_busy_s1_address),                     //                     i2c_busy_s1.address
		.i2c_busy_s1_readdata                    (mm_interconnect_0_i2c_busy_s1_readdata),                    //                                .readdata
		.i2c_dev_addr_s1_address                 (mm_interconnect_0_i2c_dev_addr_s1_address),                 //                 i2c_dev_addr_s1.address
		.i2c_dev_addr_s1_write                   (mm_interconnect_0_i2c_dev_addr_s1_write),                   //                                .write
		.i2c_dev_addr_s1_readdata                (mm_interconnect_0_i2c_dev_addr_s1_readdata),                //                                .readdata
		.i2c_dev_addr_s1_writedata               (mm_interconnect_0_i2c_dev_addr_s1_writedata),               //                                .writedata
		.i2c_dev_addr_s1_chipselect              (mm_interconnect_0_i2c_dev_addr_s1_chipselect),              //                                .chipselect
		.i2c_en_s1_address                       (mm_interconnect_0_i2c_en_s1_address),                       //                       i2c_en_s1.address
		.i2c_en_s1_write                         (mm_interconnect_0_i2c_en_s1_write),                         //                                .write
		.i2c_en_s1_readdata                      (mm_interconnect_0_i2c_en_s1_readdata),                      //                                .readdata
		.i2c_en_s1_writedata                     (mm_interconnect_0_i2c_en_s1_writedata),                     //                                .writedata
		.i2c_en_s1_chipselect                    (mm_interconnect_0_i2c_en_s1_chipselect),                    //                                .chipselect
		.i2c_miso_s1_address                     (mm_interconnect_0_i2c_miso_s1_address),                     //                     i2c_miso_s1.address
		.i2c_miso_s1_readdata                    (mm_interconnect_0_i2c_miso_s1_readdata),                    //                                .readdata
		.i2c_mosi_s1_address                     (mm_interconnect_0_i2c_mosi_s1_address),                     //                     i2c_mosi_s1.address
		.i2c_mosi_s1_write                       (mm_interconnect_0_i2c_mosi_s1_write),                       //                                .write
		.i2c_mosi_s1_readdata                    (mm_interconnect_0_i2c_mosi_s1_readdata),                    //                                .readdata
		.i2c_mosi_s1_writedata                   (mm_interconnect_0_i2c_mosi_s1_writedata),                   //                                .writedata
		.i2c_mosi_s1_chipselect                  (mm_interconnect_0_i2c_mosi_s1_chipselect),                  //                                .chipselect
		.i2c_reg_addr_s1_address                 (mm_interconnect_0_i2c_reg_addr_s1_address),                 //                 i2c_reg_addr_s1.address
		.i2c_reg_addr_s1_write                   (mm_interconnect_0_i2c_reg_addr_s1_write),                   //                                .write
		.i2c_reg_addr_s1_readdata                (mm_interconnect_0_i2c_reg_addr_s1_readdata),                //                                .readdata
		.i2c_reg_addr_s1_writedata               (mm_interconnect_0_i2c_reg_addr_s1_writedata),               //                                .writedata
		.i2c_reg_addr_s1_chipselect              (mm_interconnect_0_i2c_reg_addr_s1_chipselect),              //                                .chipselect
		.i2c_rst_s1_address                      (mm_interconnect_0_i2c_rst_s1_address),                      //                      i2c_rst_s1.address
		.i2c_rst_s1_write                        (mm_interconnect_0_i2c_rst_s1_write),                        //                                .write
		.i2c_rst_s1_readdata                     (mm_interconnect_0_i2c_rst_s1_readdata),                     //                                .readdata
		.i2c_rst_s1_writedata                    (mm_interconnect_0_i2c_rst_s1_writedata),                    //                                .writedata
		.i2c_rst_s1_chipselect                   (mm_interconnect_0_i2c_rst_s1_chipselect),                   //                                .chipselect
		.i2c_rw_s1_address                       (mm_interconnect_0_i2c_rw_s1_address),                       //                       i2c_rw_s1.address
		.i2c_rw_s1_write                         (mm_interconnect_0_i2c_rw_s1_write),                         //                                .write
		.i2c_rw_s1_readdata                      (mm_interconnect_0_i2c_rw_s1_readdata),                      //                                .readdata
		.i2c_rw_s1_writedata                     (mm_interconnect_0_i2c_rw_s1_writedata),                     //                                .writedata
		.i2c_rw_s1_chipselect                    (mm_interconnect_0_i2c_rw_s1_chipselect),                    //                                .chipselect
		.in_H_s1_address                         (mm_interconnect_0_in_h_s1_address),                         //                         in_H_s1.address
		.in_H_s1_readdata                        (mm_interconnect_0_in_h_s1_readdata),                        //                                .readdata
		.in_L_s1_address                         (mm_interconnect_0_in_l_s1_address),                         //                         in_L_s1.address
		.in_L_s1_readdata                        (mm_interconnect_0_in_l_s1_readdata),                        //                                .readdata
		.jtag_uart_avalon_jtag_slave_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //     jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write       (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),       //                                .write
		.jtag_uart_avalon_jtag_slave_read        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),        //                                .read
		.jtag_uart_avalon_jtag_slave_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                                .readdata
		.jtag_uart_avalon_jtag_slave_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                                .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                                .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  //                                .chipselect
		.led_s1_address                          (mm_interconnect_0_led_s1_address),                          //                          led_s1.address
		.led_s1_write                            (mm_interconnect_0_led_s1_write),                            //                                .write
		.led_s1_readdata                         (mm_interconnect_0_led_s1_readdata),                         //                                .readdata
		.led_s1_writedata                        (mm_interconnect_0_led_s1_writedata),                        //                                .writedata
		.led_s1_chipselect                       (mm_interconnect_0_led_s1_chipselect),                       //                                .chipselect
		.onchip_memory_s1_address                (mm_interconnect_0_onchip_memory_s1_address),                //                onchip_memory_s1.address
		.onchip_memory_s1_write                  (mm_interconnect_0_onchip_memory_s1_write),                  //                                .write
		.onchip_memory_s1_readdata               (mm_interconnect_0_onchip_memory_s1_readdata),               //                                .readdata
		.onchip_memory_s1_writedata              (mm_interconnect_0_onchip_memory_s1_writedata),              //                                .writedata
		.onchip_memory_s1_byteenable             (mm_interconnect_0_onchip_memory_s1_byteenable),             //                                .byteenable
		.onchip_memory_s1_chipselect             (mm_interconnect_0_onchip_memory_s1_chipselect),             //                                .chipselect
		.onchip_memory_s1_clken                  (mm_interconnect_0_onchip_memory_s1_clken),                  //                                .clken
		.out0_s1_address                         (mm_interconnect_0_out0_s1_address),                         //                         out0_s1.address
		.out0_s1_write                           (mm_interconnect_0_out0_s1_write),                           //                                .write
		.out0_s1_readdata                        (mm_interconnect_0_out0_s1_readdata),                        //                                .readdata
		.out0_s1_writedata                       (mm_interconnect_0_out0_s1_writedata),                       //                                .writedata
		.out0_s1_chipselect                      (mm_interconnect_0_out0_s1_chipselect),                      //                                .chipselect
		.out1_s1_address                         (mm_interconnect_0_out1_s1_address),                         //                         out1_s1.address
		.out1_s1_write                           (mm_interconnect_0_out1_s1_write),                           //                                .write
		.out1_s1_readdata                        (mm_interconnect_0_out1_s1_readdata),                        //                                .readdata
		.out1_s1_writedata                       (mm_interconnect_0_out1_s1_writedata),                       //                                .writedata
		.out1_s1_chipselect                      (mm_interconnect_0_out1_s1_chipselect),                      //                                .chipselect
		.sample_clk_s1_address                   (mm_interconnect_0_sample_clk_s1_address),                   //                   sample_clk_s1.address
		.sample_clk_s1_write                     (mm_interconnect_0_sample_clk_s1_write),                     //                                .write
		.sample_clk_s1_readdata                  (mm_interconnect_0_sample_clk_s1_readdata),                  //                                .readdata
		.sample_clk_s1_writedata                 (mm_interconnect_0_sample_clk_s1_writedata),                 //                                .writedata
		.sample_clk_s1_chipselect                (mm_interconnect_0_sample_clk_s1_chipselect)                 //                                .chipselect
	);

	unsaved_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (cpu_irq_irq)                     //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
